VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO logo
  CLASS BLOCK ;
  FOREIGN logo ;
  ORIGIN 11.960 21.580 ;
  SIZE 26.120 BY 37.500 ;
  OBS
      LAYER met5 ;
        RECT -11.960 9.350 13.000 15.920 ;
        RECT -11.680 -12.070 -5.430 5.530 ;
        RECT -0.590 -0.400 1.860 1.670 ;
        RECT -0.410 -8.590 1.840 -6.030 ;
        RECT 7.910 -11.850 14.160 5.750 ;
        RECT -11.470 -21.580 13.460 -17.470 ;
  END
END logo
END LIBRARY

