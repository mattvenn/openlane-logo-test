VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO LOGO
  CLASS BLOCK ;
  FOREIGN LOGO ;
  ORIGIN 0.000 -20.000 ;
  SIZE 800.000 BY 800.000 ;
  OBS
      LAYER met5 ;
        RECT 80.000 800.000 140.000 820.000 ;
        RECT 660.000 800.000 720.000 820.000 ;
        RECT 100.000 780.000 180.000 800.000 ;
        RECT 120.000 760.000 180.000 780.000 ;
        RECT 620.000 780.000 700.000 800.000 ;
        RECT 620.000 760.000 680.000 780.000 ;
        RECT 140.000 740.000 200.000 760.000 ;
        RECT 120.000 720.000 200.000 740.000 ;
        RECT 0.000 700.000 20.000 720.000 ;
        RECT 100.000 700.000 200.000 720.000 ;
        RECT 0.000 680.000 40.000 700.000 ;
        RECT 80.000 680.000 200.000 700.000 ;
        RECT 600.000 740.000 660.000 760.000 ;
        RECT 600.000 720.000 680.000 740.000 ;
        RECT 600.000 700.000 700.000 720.000 ;
        RECT 780.000 700.000 800.000 720.000 ;
        RECT 600.000 680.000 720.000 700.000 ;
        RECT 760.000 680.000 800.000 700.000 ;
        RECT 0.000 660.000 220.000 680.000 ;
        RECT 580.000 660.000 800.000 680.000 ;
        RECT 20.000 640.000 240.000 660.000 ;
        RECT 560.000 640.000 780.000 660.000 ;
        RECT 20.000 620.000 260.000 640.000 ;
        RECT 340.000 620.000 460.000 640.000 ;
        RECT 540.000 620.000 780.000 640.000 ;
        RECT 60.000 600.000 280.000 620.000 ;
        RECT 300.000 600.000 500.000 620.000 ;
        RECT 520.000 600.000 740.000 620.000 ;
        RECT 140.000 580.000 260.000 600.000 ;
        RECT 280.000 580.000 520.000 600.000 ;
        RECT 540.000 580.000 660.000 600.000 ;
        RECT 160.000 560.000 240.000 580.000 ;
        RECT 260.000 560.000 540.000 580.000 ;
        RECT 180.000 540.000 540.000 560.000 ;
        RECT 560.000 560.000 640.000 580.000 ;
        RECT 560.000 540.000 620.000 560.000 ;
        RECT 200.000 520.000 220.000 540.000 ;
        RECT 240.000 520.000 560.000 540.000 ;
        RECT 580.000 520.000 600.000 540.000 ;
        RECT 220.000 460.000 580.000 520.000 ;
        RECT 220.000 440.000 280.000 460.000 ;
        RECT 200.000 380.000 260.000 440.000 ;
        RECT 360.000 400.000 440.000 460.000 ;
        RECT 520.000 440.000 580.000 460.000 ;
        RECT 540.000 420.000 580.000 440.000 ;
        RECT 340.000 380.000 460.000 400.000 ;
        RECT 540.000 380.000 600.000 420.000 ;
        RECT 220.000 360.000 260.000 380.000 ;
        RECT 220.000 340.000 280.000 360.000 ;
        RECT 300.000 340.000 500.000 380.000 ;
        RECT 540.000 360.000 580.000 380.000 ;
        RECT 520.000 340.000 580.000 360.000 ;
        RECT 220.000 320.000 380.000 340.000 ;
        RECT 200.000 300.000 380.000 320.000 ;
        RECT 180.000 280.000 220.000 300.000 ;
        RECT 160.000 260.000 220.000 280.000 ;
        RECT 240.000 280.000 380.000 300.000 ;
        RECT 420.000 320.000 580.000 340.000 ;
        RECT 420.000 300.000 600.000 320.000 ;
        RECT 420.000 280.000 560.000 300.000 ;
        RECT 240.000 260.000 560.000 280.000 ;
        RECT 580.000 280.000 620.000 300.000 ;
        RECT 580.000 260.000 640.000 280.000 ;
        RECT 140.000 240.000 240.000 260.000 ;
        RECT 260.000 240.000 540.000 260.000 ;
        RECT 560.000 240.000 660.000 260.000 ;
        RECT 60.000 220.000 260.000 240.000 ;
        RECT 20.000 200.000 260.000 220.000 ;
        RECT 20.000 180.000 240.000 200.000 ;
        RECT 280.000 180.000 520.000 240.000 ;
        RECT 540.000 220.000 740.000 240.000 ;
        RECT 540.000 200.000 780.000 220.000 ;
        RECT 560.000 180.000 780.000 200.000 ;
        RECT 0.000 160.000 60.000 180.000 ;
        RECT 80.000 160.000 220.000 180.000 ;
        RECT 300.000 160.000 360.000 180.000 ;
        RECT 380.000 160.000 420.000 180.000 ;
        RECT 440.000 160.000 500.000 180.000 ;
        RECT 580.000 160.000 720.000 180.000 ;
        RECT 740.000 160.000 800.000 180.000 ;
        RECT 0.000 140.000 40.000 160.000 ;
        RECT 80.000 140.000 200.000 160.000 ;
        RECT 0.000 120.000 20.000 140.000 ;
        RECT 100.000 120.000 200.000 140.000 ;
        RECT 120.000 100.000 200.000 120.000 ;
        RECT 140.000 80.000 200.000 100.000 ;
        RECT 600.000 140.000 720.000 160.000 ;
        RECT 760.000 140.000 800.000 160.000 ;
        RECT 600.000 120.000 700.000 140.000 ;
        RECT 780.000 120.000 800.000 140.000 ;
        RECT 600.000 100.000 680.000 120.000 ;
        RECT 600.000 80.000 660.000 100.000 ;
        RECT 120.000 60.000 180.000 80.000 ;
        RECT 100.000 40.000 180.000 60.000 ;
        RECT 620.000 60.000 680.000 80.000 ;
        RECT 620.000 40.000 700.000 60.000 ;
        RECT 80.000 20.000 140.000 40.000 ;
        RECT 660.000 20.000 720.000 40.000 ;
  END
END LOGO
END LIBRARY

